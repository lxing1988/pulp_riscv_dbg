/* Copyright 2018 ETH Zurich and University of Bologna.
 * Copyright and related rights are licensed under the Solderpad Hardware
 * License, Version 0.51 (the “License”); you may not use this file except in
 * compliance with the License.  You may obtain a copy of the License at
 * http://solderpad.org/licenses/SHL-0.51. Unless required by applicable law
 * or agreed to in writing, software, hardware and materials distributed under
 * this License is distributed on an “AS IS” BASIS, WITHOUT WARRANTIES OR
 * CONDITIONS OF ANY KIND, either express or implied. See the License for the
 * specific language governing permissions and limitations under the License.
 *
 * File: $filename.v
 *
 * Description: Auto-generated 32 bits bootrom
 */

// Auto-generated code
module bootrom (
   input  logic         clk_i,
   input  logic         req_i,
   input  logic [31:0]  addr_i,
   output logic [31:0]  rdata_o
);
    localparam int RomSize = 286;

    const logic [RomSize-1:0][31:0] mem = {
        32'h00646564,
        32'h6e657478,
        32'h652d7374,
        32'h70757272,
        32'h65746e69,
        32'h00736567,
        32'h6e617200,
        32'h656c646e,
        32'h6168702c,
        32'h78756e69,
        32'h6c007265,
        32'h6c6c6f72,
        32'h746e6f63,
        32'h2d747075,
        32'h72726574,
        32'h6e690073,
        32'h6c6c6563,
        32'h2d747075,
        32'h72726574,
        32'h6e692300,
        32'h79636e65,
        32'h75716572,
        32'h662d6b63,
        32'h6f6c6300,
        32'h65707974,
        32'h2d756d6d,
        32'h00617369,
        32'h2c766373,
        32'h69720073,
        32'h75746174,
        32'h73006765,
        32'h72006570,
        32'h79745f65,
        32'h63697665,
        32'h64007963,
        32'h6e657571,
        32'h6572662d,
        32'h65736162,
        32'h656d6974,
        32'h006c6564,
        32'h6f6d0065,
        32'h6c626974,
        32'h61706d6f,
        32'h6300736c,
        32'h6c65632d,
        32'h657a6973,
        32'h2300736c,
        32'h6c65632d,
        32'h73736572,
        32'h64646123,
        32'h09000000,
        32'h02000000,
        32'h02000000,
        32'h00000030,
        32'h66697468,
        32'h2c626375,
        32'h1b000000,
        32'h0a000000,
        32'h03000000,
        32'h00000000,
        32'h66697468,
        32'h01000000,
        32'h02000000,
        32'h02000000,
        32'h00000c00,
        32'h00000000,
        32'h00000002,
        32'h00000000,
        32'h4b000000,
        32'h10000000,
        32'h03000000,
        32'h07000000,
        32'h01000000,
        32'h03000000,
        32'h01000000,
        32'hb4000000,
        32'h10000000,
        32'h03000000,
        32'h00000000,
        32'h30746e69,
        32'h6c632c76,
        32'h63736972,
        32'h1b000000,
        32'h0d000000,
        32'h03000000,
        32'h00000030,
        32'h30303030,
        32'h30324074,
        32'h6e696c63,
        32'h01000000,
        32'had000000,
        32'h00000000,
        32'h03000000,
        32'h00007375,
        32'h622d656c,
        32'h706d6973,
        32'h00636f73,
        32'h2d657261,
        32'h622d656e,
        32'h61697261,
        32'h2c687465,
        32'h1b000000,
        32'h1f000000,
        32'h03000000,
        32'h02000000,
        32'h0f000000,
        32'h04000000,
        32'h03000000,
        32'h02000000,
        32'h00000000,
        32'h04000000,
        32'h03000000,
        32'h00636f73,
        32'h01000000,
        32'h02000000,
        32'h00000001,
        32'h00000000,
        32'h00000080,
        32'h00000000,
        32'h4b000000,
        32'h10000000,
        32'h03000000,
        32'h00007972,
        32'h6f6d656d,
        32'h3f000000,
        32'h07000000,
        32'h03000000,
        32'h00303030,
        32'h30303030,
        32'h38407972,
        32'h6f6d656d,
        32'h01000000,
        32'h02000000,
        32'h02000000,
        32'h02000000,
        32'h01000000,
        32'ha5000000,
        32'h04000000,
        32'h03000000,
        32'h01000000,
        32'h9f000000,
        32'h04000000,
        32'h03000000,
        32'h00006374,
        32'h6e692d75,
        32'h70632c76,
        32'h63736972,
        32'h1b000000,
        32'h0f000000,
        32'h03000000,
        32'h8a000000,
        32'h00000000,
        32'h03000000,
        32'h01000000,
        32'h79000000,
        32'h04000000,
        32'h03000000,
        32'h00000000,
        32'h72656c6c,
        32'h6f72746e,
        32'h6f632d74,
        32'h70757272,
        32'h65746e69,
        32'h01000000,
        32'h00ca9a3b,
        32'h69000000,
        32'h04000000,
        32'h03000000,
        32'h00003933,
        32'h76732c76,
        32'h63736972,
        32'h60000000,
        32'h0b000000,
        32'h03000000,
        32'h00636d69,
        32'h34367672,
        32'h56000000,
        32'h08000000,
        32'h03000000,
        32'h00000076,
        32'h63736972,
        32'h1b000000,
        32'h06000000,
        32'h03000000,
        32'h00000000,
        32'h79616b6f,
        32'h4f000000,
        32'h05000000,
        32'h03000000,
        32'h00000000,
        32'h4b000000,
        32'h04000000,
        32'h03000000,
        32'h00757063,
        32'h3f000000,
        32'h04000000,
        32'h03000000,
        32'h00000030,
        32'h40757063,
        32'h01000000,
        32'h80969800,
        32'h2c000000,
        32'h04000000,
        32'h03000000,
        32'h00000000,
        32'h0f000000,
        32'h04000000,
        32'h03000000,
        32'h01000000,
        32'h00000000,
        32'h04000000,
        32'h03000000,
        32'h00000000,
        32'h73757063,
        32'h01000000,
        32'h00657261,
        32'h622d656e,
        32'h61697261,
        32'h2c687465,
        32'h26000000,
        32'h10000000,
        32'h03000000,
        32'h00766564,
        32'h2d657261,
        32'h622d656e,
        32'h61697261,
        32'h2c687465,
        32'h1b000000,
        32'h14000000,
        32'h03000000,
        32'h02000000,
        32'h0f000000,
        32'h04000000,
        32'h03000000,
        32'h02000000,
        32'h00000000,
        32'h04000000,
        32'h03000000,
        32'h00000000,
        32'h01000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'hf8020000,
        32'hc8000000,
        32'h00000000,
        32'h10000000,
        32'h11000000,
        32'h28000000,
        32'h30030000,
        32'h38000000,
        32'hf8030000,
        32'hedfe0dd0,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h0000bff5,
        32'h10500073,
        32'h03c58593,
        32'h00000597,
        32'hf1402573,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00000000,
        32'h00008402,
        32'h07458593,
        32'h00000597,
        32'hf1402573,
        32'h01f41413,
        32'h0010041b
    };

    logic [$clog2(RomSize)-1:0] addr_q;

    always_ff @(posedge clk_i) begin
        if (req_i) begin
            addr_q <= addr_i[$clog2(RomSize)-1+3:3];
        end
    end

    assign rdata_o = mem[addr_q];
endmodule
